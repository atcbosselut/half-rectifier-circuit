*Amplifier

*Signals
Vdd 1 0 DC 17V
*Isig 1 2 DC 1mA
Vtr 2 0 AC 1 sin(0 .05V 10000)
Cc1 2 3 4.5u

*Gate Resistances
Rg1 1 3 120k
Rg2 3 0 50k

*Drain 
Rd 1 4 26k

*Source
Rs 5 0 4600
Cs 5 0 15.7u

*NMOS
M1 4 3 5 5 nnMOS L=10u W=10u

*Load
Rl 4 0 1e6
Cl 4 0 10p

* CD4007 Discrete NMOS & PMOS
.model nnMOS NMOS (LEVEL=2 VTo=1.4 Kp=.6m LAMBDA=0.005)
.model ppMOS PMOS (LEVEL=2 VTo=-1.0 KP=.6m LAMBDA=0.01)
*Analysis Requests
*.OPTIONS ITL5 = 0
.TRAN .5ms 100ms
.AC DEC 10 .01 10Meg

.plot TRAN V(4,0)
.PROBE
.end
